module alu(A, B, ALUCtrl, Out);

	input [31:0]A;
	input [31:0]B;
	input ALUCtrl;  // operation being executed
	
	output [31:0]Out;
	
	
	
	
endmodule
