module NoiseRemove (iCLK,
					iRST,
					iBinary,
					iDVAL,
					iX_Cont, 
					iY_Cont,
					iFrame_En,
					oDCLEAN,
					oDVAL
					);

input	      	iCLK;
input			iRST;
input	    	iBinary;
input	     	iDVAL;
input	[15:0]  iX_Cont;
input	[15:0]  iY_Cont;
input			iFrame_En;
output 	    	oDCLEAN;
output			oDVAL;

// code starts from here

endmodule