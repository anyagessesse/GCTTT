module MovementDetection (iCLK,
					      iRST,
					      iDVAL,
					      iFT_X,
					      iFT_Y, 
					      iFrame_En,
					      oGrid_Num,
					      oStable_hand,
					      );

input	      	iCLK;
input			iRST;
input	     	iDVAL;
input	[9:0]   iFT_X;
input	[9:0]   iFT_Y;
input			iFrame_En;
output 	[3:0]   oGrid_Num;
output			oStable_hand;

// code starts from here

endmodule