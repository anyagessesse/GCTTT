module Source2Binary (iCLK,
					iRST,
					iDATA,
					iDVAL,
					iX_Cont, 
					iY_Cont,
					iFrame_En,
					oBinary,
					oDVAL
					);

input	      	iCLK;
input			iRST;
input	[11:0]	iDATA;
input	     	iDVAL;
input	[15:0]  iX_Cont;
input	[15:0]  iY_Cont;
input			iFrame_En;
output 	    	oBinary;
output			oDVAL;

// code starts from here

endmodule