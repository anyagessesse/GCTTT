module FrameCapture (iCLK,
					iRST,
					iFVAL,
					oFrame_En,
					);

input	      	iCLK;
input			iRST;
input			iFVAL;
output			oFrame_En;

// code starts here

endmodule