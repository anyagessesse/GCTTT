module jumpbranch();

	input EQ;
	input LT;
	input GT;
	input LE;
	input GE;
	input NE;
	input JumpOrBranchHigh;
	input instr;
	
	output SelectJOrB;
	output flush;
	
	// decide if we should branch based on opcode & condition codes
	




endmodule

